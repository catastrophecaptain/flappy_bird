`timescale 1ps / 1ps
module control (
    input wire clk,  //时钟
    input wire rst,  //rst为1时游戏重新开始
    input up,  //up为1时小鸟飞起，连接btn
    //input mode,  //mode为1时双人模式，为0时单人模式
    input pipe_up,
    input pipe_down,
    output reg [1:0]status,  
    output reg [15:0]score,  //分数
    output reg [15:0]bird_y, //bird_y为小鸟下侧y坐标，第16位记录小鸟是否在下落，为0时小鸟下落，为1时小鸟上升
    output reg [31:0]pipe1,//pipe1储存管道1的x和y和gap，x占高10位，y占低10位，x为管子左边界坐标，y为管子上侧坐标
    output reg [31:0]pipe2,//pipe2储存管道2的x和y和gap，x占高10位，y占低10位，x为管子左边界坐标，y为管子上侧坐标
    output reg [31:0]pipe3,//pipe3储存管道3的x和y和gap，x占高10位，y占低10位，x为管子左边界坐标，y为管子上侧坐标
    output reg [31:0]coin//coin储存金币的x和y，y占高10位，x占低10位，x为金币左边界坐标，y为金币下侧坐标
	 //output reg [3:0]bird_falling
);
  wire [31:0] clk_div;
  // wire up1;
  // wire pipeup1;
  // wire pipedown1;
  reg [1:0]cnt=3;
  reg fail;//fail为1游戏结束
  //reg pass1;
  //reg pass2;
  //reg pass3; //pass1,pass2,pass3为小鸟是否通过管道，为1时通过
  reg longpress;
  reg [9:0] pipe1_x;  //pipe1_x为管1的x左边界坐标
  reg [9:0] pipe1_y;  //pipe1_y为管1的y上边界坐标
  reg [9:0] pipe2_x;  //pipe2_x为管2的x左边界坐标
  reg [9:0] pipe2_y;  //pipe2_y为管2的y上边界坐标
  reg [9:0] pipe3_x;  //pipe3_x为管3的x左边界坐标
  reg [9:0] pipe3_y;  //pipe3_y为管3的y上边界坐标
  wire [9:0] bird_x = 10'd70;  //bird_x为小鸟左边界坐标，小鸟是不动的，所以x坐标为常数
  //wire [9:0] gap = 10'd50;  //gap为管道间隙，供小鸟通过
  wire [9:0] bird_width = 10'd16;  //bird_width为小鸟宽度
  wire [9:0] bird_height = 10'd16;  //bird_height为小鸟高度
  wire [9:0] pipe_width = 10'd50;  //pipe_width为管道宽度
  wire [7:0] pipe_head=8'd40;
  wire [7:0] coin_length=8'd16;
  reg [7:0]gap1;  //gap1为管道1的间隙，供小鸟通过
  reg [7:0]gap2;  //gap2为管道2的间隙，供小鸟通过
  reg [7:0]gap3;  //gap3为管道3的间隙，供小鸟通过
  reg [15:0] bird_flying;  //bird_flying为小鸟距离开始下落的时间，为0时小鸟下落
  reg old;
  wire clk_100ms;
  //reg bird_falltime;

  clk_div m0 (
      .clk(clk),
      .rst(1'b0),
      .clk_div(clk_div)
  );  //时钟分频，将时钟分频100ms
  // pbdebounce m1 (
  //     .clk_1ms(clk_div[17]),
  //     .btn(up),
  //     .pbreg(up1)
  // );  //按钮去抖动，将按钮信号去抖动
  // pbdebounce m3 (
  //     .clk_1ms(clk_div[17]),
  //     .btn(pipe_up),
  //     .pbreg(pipeup1)
  // );  //按钮去抖动，将按钮信号去抖动
  // pbdebounce m4 (
  //     .clk_1ms(clk_div[17]),
  //     .btn(pipe_down),
  //     .pbreg(pipedown1)
  // );  //按钮去抖动，将按钮信号去抖动
  clk_100ms m2 (
      .clk(clk),
      .clk_100ms(clk_100ms)
  );  //100ms时钟
  initial begin
    status <= 2'b01;
  end
  always @(posedge clk_100ms) begin
    if (!rst) begin
      if(status==0||status==3)status<=1;
      if(pipe_up||pipe_down) begin
        if(old==0)begin
          if(status==1)status <= 2'b10;
          else status <= 2'b01;
        end
        old <= 1;
      end
      else old <= 0;
      bird_y[14:0] <= 16'd240;  //小鸟初始位置
      bird_y[15] <= 1'b0;
      pipe1_x <= 20'd210;
      pipe2_x <= 20'd420;
      pipe3_x <= 20'd630;
      cnt <= 3;
      //pass1 <= 0;
      //pass2 <= 0;
      //pass3 <= 0;//pass1,pass2,pass3为小鸟是否通过管道，为1时通过
      //bird_falltime <= 0;
      longpress <= 0;
      fail <= 0;
      score <= 16'd0;
      bird_flying <= 16'b0000;  //小鸟距离开始下落的时间，为0时小鸟下落
      coin[31] <= 1'b1;
      coin[9:0] <= 10'd650+pipe_width+clk_div % 20;
      coin[19:10] <= 20+(clk_div+50)%(440-coin_length);
      pipe1_y <= pipe_head + clk_div % (310-pipe_head-pipe_head);  // 生成pipe_head到480-150-pipe_head的随机数
      pipe2_y <= pipe_head + (clk_div+10) % (310-pipe_head-pipe_head);  // 生成pipe_head到480-150-pipe_head的随机数
      pipe3_y <= pipe_head + (clk_div+20) % (310-pipe_head-pipe_head);  // 生成pipe_head到480-150-pipe_head的随机数
      gap1 <= 100 + clk_div % 50;
      gap2 <= 100 + (clk_div+10) % 50;
      gap3 <= 100 + (clk_div+20) % 50;
      pipe1 <= {gap1,pipe1_x, pipe1_y};
      pipe2 <= {gap2,pipe2_x, pipe2_y};
      pipe3 <= {gap3,pipe3_x, pipe3_y};
    end else begin
      if(status==1)status <= 2'b00;
      if(status==2)status <= 2'b11;
      if  (pipe_up&&!fail&&status==3)begin
        case(cnt)
          1:if(pipe1_y>=pipe_head)pipe1_y<=pipe1_y-1;
          2:if(pipe2_y>=pipe_head)pipe2_y<=pipe2_y-1;
          3:if(pipe3_y>=pipe_head)pipe3_y<=pipe3_y-1;
        endcase
      end
      if (pipe_down&&!fail&&status==3)begin
        case(cnt)
          1:if(pipe1_y+pipe_head<=330)pipe1_y<=pipe1_y+1;
          2:if(pipe2_y+pipe_head<=330)pipe2_y<=pipe2_y+1;
          3:if(pipe3_y+pipe_head<=330)pipe3_y<=pipe3_y+1;
        endcase
      end
      if (up && !fail &&!longpress) begin  //按钮按下时up为1，小鸟飞行4个周期
        bird_flying <= 16'd10;
        bird_y[15]   <= 1'b1;
        longpress <= 1;
        //bird_falltime <= 0;
      end
      if ((bird_flying<=0)||fail) begin  //小鸟下落
        bird_y[14:0] <= bird_y[14:0] + 4;
        bird_y[15] <= 1'b0;
        //bird_falltime <= bird_falltime + 1;
      end
      if ((bird_flying>0)&&(!fail)) begin  //小鸟按惯性向上飞
        bird_y[14:0] <= bird_y[14:0] - bird_flying;
        bird_flying <= bird_flying - 1;
        bird_y[15] <= 1'b1;
      end
      if (!up) begin
        longpress <= 0;
      end
      if (!fail) begin  //若游戏未结束，管道移动
        pipe1_x <= pipe1_x - 2;
        pipe2_x <= pipe2_x - 2;
        pipe3_x <= pipe3_x - 2;
        coin[9:0] <= coin[9:0] - 2;
      end
      if (pipe1_x<= 2) begin  //管道移出屏幕后重新生成
        pipe1_x <= 20'd640;
        pipe1_y <= pipe_head + clk_div % (310-pipe_head-pipe_head);  // 生成pipe_head到480-150-pipe_head的随机数
        gap1 <= 120 + clk_div % 50;
        //pass1 <= 0;
        cnt <= 1;
      end
      if (pipe2_x<= 2) begin  //管道移出屏幕后重新生成 
        pipe2_x <= 20'd640;
        pipe2_y <= pipe_head + clk_div % (310-pipe_head-pipe_head);  // 生成pipe_head到480-150-pipe_head的随机数
        gap2 <= 120 + clk_div % 50;
        //pass2 <= 0;
        cnt <= 2;
      end
      if (pipe3_x<= 2) begin  //管道移出屏幕后重新生成
        pipe3_x <= 20'd640;
        pipe3_y <= pipe_head + clk_div % (310-pipe_head-pipe_head);  // 生成pipe_head到480-150-pipe_head的随机数
        gap3 <= 120 + clk_div % 50;
        //pass3 <= 0;
        cnt <= 3;
      end
      if(coin[31]==0||coin[9:0]<=0) begin
        coin[31] <= 1'b1;
        case(cnt)
          1:coin[9:0] <= pipe1_x+pipe_width+clk_div % 20;
          2:coin[9:0] <= pipe2_x+pipe_width+clk_div % 20;
          3:coin[9:0] <= pipe3_x+pipe_width+clk_div % 20;
        endcase 
        coin[19:10] <= 20+(clk_div+50)%(440-coin_length);
      end
      if ((((bird_y[14:0] <= pipe1_y)||(bird_y[14:0]+bird_height>=pipe1_y+gap1))&&(bird_x<=pipe1_x+pipe_width)&&(bird_x+bird_width>=pipe1_x))
                ||(((bird_y[14:0] <= pipe2_y)||(bird_y[14:0]+bird_height>=pipe2_y+gap2))&&(bird_x<=pipe2_x+pipe_width)&&(bird_x+bird_width>=pipe2_x))
                ||(((bird_y[14:0] <= pipe3_y)||(bird_y[14:0]+bird_height>=pipe3_y+gap3))&&(bird_x<=pipe3_x+pipe_width)&&(bird_x+bird_width>=pipe3_x))) begin
        //若小鸟与管道相撞，游戏结束
        fail <= 1;
      end
      if (!fail) begin
        if(bird_x==pipe1_x+pipe_width) begin
          score <= score + 1;
          //pass1 <= 1;
        end
        if(bird_x==pipe2_x+pipe_width) begin
          score <= score + 1;
          //pass2 <= 1;
        end
        if(bird_x==pipe3_x+pipe_width) begin
          score <= score + 1;
          //pass3 <= 1;
        end
        //若小鸟通过管道，分数加1
      end
      if(coin[31]&&((bird_y[14:0]<=coin[19:10]+coin_length)&&(bird_y[14:0]+bird_height>=coin[19:10])&&(bird_x<=coin[9:0]+coin_length)&&(bird_x+bird_width>=coin[9:0]))) begin
        coin[31] <= 1'b0;
        score <= score + 2;
      end
      pipe1 <= {gap1,pipe1_x, pipe1_y};
      pipe2 <= {gap2,pipe2_x, pipe2_y};
      pipe3 <= {gap3,pipe3_x, pipe3_y};
    end
  end
endmodule
