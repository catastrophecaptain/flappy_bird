module keyboard (
    input wire clk,
    input wire kb_clk,
    input wire data,
    output wire [7:0] keycode,
    output wire sign
);
endmodule
